module seven_segment(
	input wire[3:0]i,
	output reg[6:0]o
);

// HEX out - rewire DE1
//  ---0---
// |       |
// 5       1
// |       |
//  ---6---
// |       |
// 4       2
// |       |
//  ---3---
always @ (*) begin
	i = i/3;
	case(i)
	
		4'b0000: o = 7'b1000000;
		4'b0001: o = 7'b1111001; //1001111
		4'b0010: o = 7'b0100100; //0010010
		4'b0011: o = 7'b0110000; //0000110
		4'b0100: o = 7'b0011001; //1001100
		4'b0101: o = 7'b0010010; //0100100
		4'b0110: o = 7'b0000010; //0100000
		4'b0111: o = 7'b1111000; //0001111
		4'b1000: o = 7'b0000000;
		4'b1001: o = 7'b0011000; //0001100
		4'b1010: o = 7'b0001000;
		4'b1011: o = 7'b0000011; //1100000
		4'b1100: o = 7'b1000110; //0110001
		4'b1101: o = 7'b0100001; //1000010
		4'b1110: o = 7'b0000110; //0110000
		4'b1111: o = 7'b0001110; //0111000
		
		//default: HEX0 = 7'b0000001;
		
		endcase
		end
		


endmodule